module essai();

initial
    begin
        $display("Debut de la simulation");
    
        $finish;
    end

endmodule
